module sub4 (s,a,b);
output [4:0] s;
input [3:0] a,b;
assign s = a-b;
endmodule
